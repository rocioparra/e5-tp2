-- Copyright (C) 2019  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 19.1.0 Build 670 09/22/2019 SJ Lite Edition"
-- CREATED		"Sat Jun 06 13:47:12 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY MUX_11b IS 
	PORT
	(
		SEL :  IN  STD_LOGIC;
		INA :  IN  STD_LOGIC_VECTOR(10 DOWNTO 0);
		INB :  IN  STD_LOGIC_VECTOR(10 DOWNTO 0);
		ADDR_OUT :  OUT  STD_LOGIC_VECTOR(10 DOWNTO 0)
	);
END MUX_11b;

ARCHITECTURE bdf_type OF MUX_11b IS 

SIGNAL	ADDR_OUT_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_9 <= INA(4) AND SEL;


SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_33 AND INB(4);


SYNTHESIZED_WIRE_29 <= INA(2) AND SEL;


SYNTHESIZED_WIRE_32 <= INA(1) AND SEL;


SYNTHESIZED_WIRE_3 <= INA(0) AND SEL;


SYNTHESIZED_WIRE_2 <= SYNTHESIZED_WIRE_33 AND INB(0);


ADDR_OUT_ALTERA_SYNTHESIZED(0) <= SYNTHESIZED_WIRE_2 OR SYNTHESIZED_WIRE_3;


SYNTHESIZED_WIRE_6 <= INA(5) AND SEL;


SYNTHESIZED_WIRE_5 <= SYNTHESIZED_WIRE_33 AND INB(5);


ADDR_OUT_ALTERA_SYNTHESIZED(5) <= SYNTHESIZED_WIRE_5 OR SYNTHESIZED_WIRE_6;


SYNTHESIZED_WIRE_11 <= INA(6) AND SEL;


SYNTHESIZED_WIRE_10 <= SYNTHESIZED_WIRE_33 AND INB(6);


ADDR_OUT_ALTERA_SYNTHESIZED(4) <= SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9;


ADDR_OUT_ALTERA_SYNTHESIZED(6) <= SYNTHESIZED_WIRE_10 OR SYNTHESIZED_WIRE_11;


SYNTHESIZED_WIRE_14 <= INA(7) AND SEL;


SYNTHESIZED_WIRE_13 <= SYNTHESIZED_WIRE_33 AND INB(7);


ADDR_OUT_ALTERA_SYNTHESIZED(7) <= SYNTHESIZED_WIRE_13 OR SYNTHESIZED_WIRE_14;


SYNTHESIZED_WIRE_17 <= INA(8) AND SEL;


SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_33 AND INB(8);


ADDR_OUT_ALTERA_SYNTHESIZED(8) <= SYNTHESIZED_WIRE_16 OR SYNTHESIZED_WIRE_17;


SYNTHESIZED_WIRE_20 <= INA(9) AND SEL;


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_33 AND INB(9);


ADDR_OUT_ALTERA_SYNTHESIZED(9) <= SYNTHESIZED_WIRE_19 OR SYNTHESIZED_WIRE_20;


SYNTHESIZED_WIRE_26 <= INA(3) AND SEL;


SYNTHESIZED_WIRE_23 <= INA(10) AND SEL;


SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_33 AND INB(10);


ADDR_OUT_ALTERA_SYNTHESIZED(10) <= SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_23;


SYNTHESIZED_WIRE_33 <= NOT(SEL);



SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_33 AND INB(3);


ADDR_OUT_ALTERA_SYNTHESIZED(3) <= SYNTHESIZED_WIRE_25 OR SYNTHESIZED_WIRE_26;


SYNTHESIZED_WIRE_28 <= SYNTHESIZED_WIRE_33 AND INB(2);


ADDR_OUT_ALTERA_SYNTHESIZED(2) <= SYNTHESIZED_WIRE_28 OR SYNTHESIZED_WIRE_29;


SYNTHESIZED_WIRE_31 <= SYNTHESIZED_WIRE_33 AND INB(1);


ADDR_OUT_ALTERA_SYNTHESIZED(1) <= SYNTHESIZED_WIRE_31 OR SYNTHESIZED_WIRE_32;

ADDR_OUT <= ADDR_OUT_ALTERA_SYNTHESIZED;

END bdf_type;