LIBRARY IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;   -- Needed for shifts

ENTITY CheckBraRet IS 
    PORT
    (
			instr_id    :  IN  STD_LOGIC_VECTOR(6 downto 0);
			BRA    		:  OUT STD_LOGIC:= '0';
			RET    		:  OUT STD_LOGIC:= '0'
    );
END CheckBraRet;

ARCHITECTURE behaviour OF CheckBraRet IS    
begin
	BRA <= '1' when(instr_id(6 downto 3) = "0111") else '0';		--BSR
	RET <= '1' when(instr_id(6 downto 0) = "0000011") else '0'; 	--RTI
END behaviour;